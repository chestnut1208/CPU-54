`timescale 1ns / 1ps

module MULTU(
    //input clk,
   // input reset,
    input [31:0] a,//multiplicand������
    input [31:0] b,//multiplier����
    output [63:0] z
    );
    
  // wire [63:0] a_ext;
   reg [63:0] mid [31:0]; //32���ӷ�����Ĵ���
   reg [63:0] add1 [15:0]; //add01�Ĵ���
   reg [63:0] add2 [7:0];
   reg [63:0] add3 [3:0];
   reg [63:0] add4 [1:0];
   reg [63:0] temp;
  // assign a_ext={32'd0,a};
   
   always@(*)
   begin
   //reset�͵�ƽ��Ч
  /* if(!reset) begin
       mid[0]<=0;
       mid[1]<=0;
       mid[2]<=0;
       mid[3]<=0;
       mid[4]<=0;
       mid[5]<=0;
       mid[6]<=0;
       mid[7]<=0;
       mid[8]<=0;
       mid[9]<=0;
       mid[10]<=0;
       mid[11]<=0;
       mid[12]<=0;
       mid[13]<=0;
       mid[14]<=0;
       mid[15]<=0;
       mid[16]<=0;
       mid[17]<=0;
       mid[18]<=0;
       mid[19]<=0;
       mid[20]<=0;
       mid[21]<=0;
       mid[22]<=0;
       mid[23]<=0;
       mid[24]<=0;
       mid[25]<=0;
       mid[26]<=0;
       mid[27]<=0;
       mid[28]<=0;
       mid[29]<=0;
       mid[30]<=0;
       mid[31]<=0;
       temp<=0;
   end
   else begin//reset�ߵ�ƽ*/
       mid[0]<=a&{(2*32){b[0]}}; //����32���ӷ�����
       mid[1]<=(a<<1) & {(2*32){b[1]}};//����b[i]��ֵ0/1�����и�ֵ+��λ
       mid[2]<=(a<<2) & {(2*32){b[2]}};
       mid[3]<=(a<<3) & {(2*32){b[3]}};
       mid[4]<=(a<<4) & {(2*32){b[4]}};
       mid[5]<=(a<<5) & {(2*32){b[5]}};
       mid[6]<=(a<<6) & {(2*32){b[6]}};
       mid[7]<=(a<<7) & {(2*32){b[7]}};
       mid[8]<=(a<<8) & {(2*32){b[8]}};
       mid[9]<=(a<<9) & {(2*32){b[9]}};
       mid[10]<=(a<<10) & {(2*32){b[10]}};
       mid[11]<=(a<<11) & {(2*32){b[11]}};
       mid[12]<=(a<<12) & {(2*32){b[12]}};
       mid[13]<=(a<<13) & {(2*32){b[13]}};
       mid[14]<=(a<<14) & {(2*32){b[14]}};
       mid[15]<=(a<<15) & {(2*32){b[15]}};
       mid[16]<=(a<<16) & {(2*32){b[16]}};
       mid[17]<=(a<<17) & {(2*32){b[17]}};
       mid[18]<=(a<<18) & {(2*32){b[18]}};
       mid[19]<=(a<<19) & {(2*32){b[19]}};
       mid[20]<=(a<<20) & {(2*32){b[20]}};
       mid[21]<=(a<<21) & {(2*32){b[21]}};
       mid[22]<=(a<<22) & {(2*32){b[22]}};
       mid[23]<=(a<<23) & {(2*32){b[23]}};
       mid[24]<=(a<<24) & {(2*32){b[24]}};
       mid[25]<=(a<<25) & {(2*32){b[25]}};
       mid[26]<=(a<<26) & {(2*32){b[26]}};
       mid[27]<=(a<<27) & {(2*32){b[27]}};
       mid[28]<=(a<<28) & {(2*32){b[28]}};
       mid[29]<=(a<<29) & {(2*32){b[29]}};
       mid[30]<=(a<<30) & {(2*32){b[30]}};
       mid[31]<=(a<<31) & {(2*32){b[31]}};
       
       add1[0]<=mid[0]+mid[1];
       add1[1]<=mid[2]+mid[3];
       add1[2]<=mid[4]+mid[5];
       add1[3]<=mid[6]+mid[7];
       add1[4]<=mid[8]+mid[9];
       add1[5]<=mid[10]+mid[11];
       add1[6]<=mid[12]+mid[13];
       add1[7]<=mid[14]+mid[15];
       add1[8]<=mid[16]+mid[17];
       add1[9]<=mid[18]+mid[19];
       add1[10]<=mid[20]+mid[21];
       add1[11]<=mid[22]+mid[23];
       add1[12]<=mid[24]+mid[25];
       add1[13]<=mid[26]+mid[27];
       add1[14]<=mid[28]+mid[29];
       add1[15]<=mid[30]+mid[31];
       
       add2[0]<=add1[0]+add1[1];
       add2[1]<=add1[2]+add1[3];
       add2[2]<=add1[4]+add1[5];
       add2[3]<=add1[6]+add1[7];
       add2[4]<=add1[8]+add1[9];
       add2[5]<=add1[10]+add1[11];
       add2[6]<=add1[12]+add1[13];
       add2[7]<=add1[14]+add1[15];
       
       add3[0]<=add2[0]+add2[1];
       add3[1]<=add2[2]+add2[3];
       add3[2]<=add2[4]+add2[5];
       add3[3]<=add2[6]+add2[7];
       
       add4[0]<=add3[0]+add3[1];
       add4[1]<=add3[2]+add3[3];
       
       temp<=add4[0]+add4[1];
       
   end//end of else
   //end//end of always
   assign z=temp;
   
endmodule
